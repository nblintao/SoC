// data length is 128
// ram depth is 7
module mio_rom (a, inst, rom_a, d_f_rom);
    input  [31:0] a;
    output [31:0] inst; 
    input  [31:0] rom_a;
    output [31:0] d_f_rom;

    wire   [31:0] rom [0:127];
    assign inst    = rom[a[8:2]];
    assign d_f_rom = rom[rom_a[8:2]];

    assign rom[7'h00] = 32'b00100000000111010001000000000000;
    assign rom[7'h01] = 32'b00100011101111011111111111101100;
    assign rom[7'h02] = 32'b10101111101000000000000000000000;
    assign rom[7'h03] = 32'b10101111101000000000000000000100;
    assign rom[7'h04] = 32'b00100000000010000000000000110010;
    assign rom[7'h05] = 32'b10101111101010000000000000001000;
    assign rom[7'h06] = 32'b10101111101010000000000000001100;
    assign rom[7'h07] = 32'b00100000000010000000000000000001;
    assign rom[7'h08] = 32'b10101111101010000000000000010000;
    assign rom[7'h09] = 32'b00100000000010000000000000011111;
    assign rom[7'h0a] = 32'b00111100000010011100000000000000;
    assign rom[7'h0b] = 32'b00110101001010010000000000000000;
    assign rom[7'h0c] = 32'b10101101001010000000000000000000;
    assign rom[7'h0d] = 32'b00000000000111010010100000100000;
    assign rom[7'h0e] = 32'b00111100000010001010000000000000;
    assign rom[7'h0f] = 32'b00110101000010000000000000000000;
    assign rom[7'h10] = 32'b10001101000100000000000000000000;
    assign rom[7'h11] = 32'b00110010000010000000000100000000;
    assign rom[7'h12] = 32'b00010001000000000000000000000010;
    assign rom[7'h13] = 32'b00000000000100000010000000000000;
    assign rom[7'h14] = 32'b00001100000000000000000001000001;
    assign rom[7'h15] = 32'b10001100000010000001000000001000;
    assign rom[7'h16] = 32'b00010101000000000000000000000001;
    assign rom[7'h17] = 32'b00001100000000000000000000011001;
    assign rom[7'h18] = 32'b00001000000000000000000000001101;
    assign rom[7'h19] = 32'b10001100101010000000000000001100;
    assign rom[7'h1a] = 32'b00010001000000000000000000000011;
    assign rom[7'h1b] = 32'b00100001000010001111111111111111;
    assign rom[7'h1c] = 32'b10101100101010000000000000001100;
    assign rom[7'h1d] = 32'b00000011111000000000000000001000;
    assign rom[7'h1e] = 32'b10001100101010000000000000001000;
    assign rom[7'h1f] = 32'b10101100101010000000000000001100;
    assign rom[7'h20] = 32'b10001100101010100000000000000000;
    assign rom[7'h21] = 32'b10001100101010110000000000000100;
    assign rom[7'h22] = 32'b10001100101011000000000000010000;
    assign rom[7'h23] = 32'b00100000000010010000000001001111;
    assign rom[7'h24] = 32'b00010101001010110000000000000011;
    assign rom[7'h25] = 32'b00000000000011000100100000101010;
    assign rom[7'h26] = 32'b00010001001000000000000000000001;
    assign rom[7'h27] = 32'b00001000000000000000000000101100;
    assign rom[7'h28] = 32'b00100000000010010000000000000000;
    assign rom[7'h29] = 32'b00010101001010110000000000000101;
    assign rom[7'h2a] = 32'b00000001100000000100100000101010;
    assign rom[7'h2b] = 32'b00010001001000000000000000000011;
    assign rom[7'h2c] = 32'b00000000000011000110000000100010;
    assign rom[7'h2d] = 32'b10101100101011000000000000001000;
    assign rom[7'h2e] = 32'b00001000000000000000000001000000;
    assign rom[7'h2f] = 32'b00100011101111011111111111110100;
    assign rom[7'h30] = 32'b10101111101001000000000000000000;
    assign rom[7'h31] = 32'b10101111101001010000000000000100;
    assign rom[7'h32] = 32'b10101111101111110000000000001000;
    assign rom[7'h33] = 32'b00000000000010100010000000000000;
    assign rom[7'h34] = 32'b00000000000010110010100000000000;
    assign rom[7'h35] = 32'b00000000000011000110100000101010;
    assign rom[7'h36] = 32'b00010001101000000000000000000010;
    assign rom[7'h37] = 32'b00001100000000000000000001100000;
    assign rom[7'h38] = 32'b00001000000000000000000000111010;
    assign rom[7'h39] = 32'b00001100000000000000000001101111;
    assign rom[7'h3a] = 32'b10001111101001000000000000000000;
    assign rom[7'h3b] = 32'b10001111101001010000000000000100;
    assign rom[7'h3c] = 32'b10001111101111110000000000001000;
    assign rom[7'h3d] = 32'b00100011101111010000000000001100;
    assign rom[7'h3e] = 32'b10101100101000100000000000000000;
    assign rom[7'h3f] = 32'b10101100101000110000000000000100;
    assign rom[7'h40] = 32'b00000011111000000000000000001000;
    assign rom[7'h41] = 32'b00100011101111011111111111111100;
    assign rom[7'h42] = 32'b10101111101111110000000000000000;
    assign rom[7'h43] = 32'b00100000000010000001000000000010;
    assign rom[7'h44] = 32'b10001101000010010000000000000000;
    assign rom[7'h45] = 32'b00010101001000000000000000010110;
    assign rom[7'h46] = 32'b00111100000010010000000000000000;
    assign rom[7'h47] = 32'b00110101001010010000000111110000;
    assign rom[7'h48] = 32'b00010001001001000000000000010001;
    assign rom[7'h49] = 32'b00110000100001000000000011111111;
    assign rom[7'h4a] = 32'b00100000000010100000000001110100;
    assign rom[7'h4b] = 32'b00010001010001000000000000000001;
    assign rom[7'h4c] = 32'b00001000000000000000000001011101;
    assign rom[7'h4d] = 32'b00100011101111011111111111111000;
    assign rom[7'h4e] = 32'b10101111101001000000000000000000;
    assign rom[7'h4f] = 32'b10101111101001010000000000000100;
    assign rom[7'h50] = 32'b00000000000001010100000000000000;
    assign rom[7'h51] = 32'b10001101000001000000000000000000;
    assign rom[7'h52] = 32'b10001101000001010000000000000100;
    assign rom[7'h53] = 32'b00001100000000000000000001100000;
    assign rom[7'h54] = 32'b10001111101001000000000000000000;
    assign rom[7'h55] = 32'b10001111101001010000000000000100;
    assign rom[7'h56] = 32'b00100011101111010000000000001000;
    assign rom[7'h57] = 32'b10101100101000100000000000000000;
    assign rom[7'h58] = 32'b10101100101000110000000000000100;
    assign rom[7'h59] = 32'b00001000000000000000000001011101;
    assign rom[7'h5a] = 32'b10101101000010010000000000000000;
    assign rom[7'h5b] = 32'b00001000000000000000000001011101;
    assign rom[7'h5c] = 32'b10101101000000000000000000000000;
    assign rom[7'h5d] = 32'b10001111101111110000000000000000;
    assign rom[7'h5e] = 32'b00100011101111010000000000000100;
    assign rom[7'h5f] = 32'b00000011111000000000000000001000;
    assign rom[7'h60] = 32'b00000000000001000100000110000000;
    assign rom[7'h61] = 32'b00000000000001000100100100000000;
    assign rom[7'h62] = 32'b00000001000010010100000000100000;
    assign rom[7'h63] = 32'b00000001000001010100000000100000;
    assign rom[7'h64] = 32'b00000000000010000100000010000000;
    assign rom[7'h65] = 32'b00111100000010011100000000000000;
    assign rom[7'h66] = 32'b00110101001010010000000000000000;
    assign rom[7'h67] = 32'b00000001001010000100100000100000;
    assign rom[7'h68] = 32'b10001101001010100000000000000000;
    assign rom[7'h69] = 32'b10101101001000000000000000000000;
    assign rom[7'h6a] = 32'b00100000100000100000000000000000;
    assign rom[7'h6b] = 32'b00100000101000110000000000000001;
    assign rom[7'h6c] = 32'b00100001001010010000000000000100;
    assign rom[7'h6d] = 32'b10101101001010100000000000000000;
    assign rom[7'h6e] = 32'b00000011111000000000000000001000;
    assign rom[7'h6f] = 32'b00000000000001000100000110000000;
    assign rom[7'h70] = 32'b00000000000001000100100100000000;
    assign rom[7'h71] = 32'b00000001000010010100000000100000;
    assign rom[7'h72] = 32'b00000001000001010100000000100000;
    assign rom[7'h73] = 32'b00000000000010000100000010000000;
    assign rom[7'h74] = 32'b00111100000010011100000000000000;
    assign rom[7'h75] = 32'b00110101001010010000000000000000;
    assign rom[7'h76] = 32'b00000001001010000100100000100000;
    assign rom[7'h77] = 32'b10001101001010100000000000000000;
    assign rom[7'h78] = 32'b10101101001000000000000000000000;
    assign rom[7'h79] = 32'b00100000100000100000000000000000;
    assign rom[7'h7a] = 32'b00100000101000111111111111111111;
    assign rom[7'h7b] = 32'b00100001001010011111111111111100;
    assign rom[7'h7c] = 32'b10101101001010100000000000000000;
    assign rom[7'h7d] = 32'b00000011111000000000000000001000;
    assign rom[7'h7e] = 32'b00001000000000000000000001111110;
    assign rom[7'h7f] = 32'b00000000000000000000000000000000;
endmodule
