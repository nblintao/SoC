module inst_mem_v (a,inst);   // instruction memory, rom
    input  [31:0] a;                        // address
    output [31:0] inst;                     // instruction
    wire   [31:0] rom [0:63];               // rom cells: 64 words * 32 bits
    assign inst = rom[a[7:2]];              // use word address to read rom
    // rom[word_addr] = instruction
assign rom[6'h0] = 32'b00111100000000111100000000000000;
assign rom[6'h1] = 32'b00100000000001010000000000100001;
assign rom[6'h2] = 32'b00001100000000000000000000000111;
assign rom[6'h3] = 32'b00100000101001010000000000000001;
assign rom[6'h4] = 32'b00101000101000100000000000101000;
assign rom[6'h5] = 32'b00010100010000001111111111111100;
assign rom[6'h6] = 32'b00001000000000000000000000000110;
assign rom[6'h7] = 32'b10101100011001010000000000000000;
assign rom[6'h8] = 32'b00100000011000110000000000000100;
assign rom[6'h9] = 32'b00000011111000000000000000001000;
assign rom[6'ha] = 32'b00000000000000000000000000000000;
assign rom[6'hb] = 32'b00000000000000000000000000000000;
assign rom[6'hc] = 32'b00000000000000000000000000000000;
assign rom[6'hd] = 32'b00000000000000000000000000000000;
assign rom[6'he] = 32'b00000000000000000000000000000000;
assign rom[6'hf] = 32'b00000000000000000000000000000000;
assign rom[6'h10] = 32'b00000000000000000000000000000000;
assign rom[6'h11] = 32'b00000000000000000000000000000000;
assign rom[6'h12] = 32'b00000000000000000000000000000000;
assign rom[6'h13] = 32'b00000000000000000000000000000000;
assign rom[6'h14] = 32'b00000000000000000000000000000000;
assign rom[6'h15] = 32'b00000000000000000000000000000000;
assign rom[6'h16] = 32'b00000000000000000000000000000000;
assign rom[6'h17] = 32'b00000000000000000000000000000000;
assign rom[6'h18] = 32'b00000000000000000000000000000000;
assign rom[6'h19] = 32'b00000000000000000000000000000000;
assign rom[6'h1a] = 32'b00000000000000000000000000000000;
assign rom[6'h1b] = 32'b00000000000000000000000000000000;
assign rom[6'h1c] = 32'b00000000000000000000000000000000;
assign rom[6'h1d] = 32'b00000000000000000000000000000000;
assign rom[6'h1e] = 32'b00000000000000000000000000000000;
assign rom[6'h1f] = 32'b00000000000000000000000000000000;
assign rom[6'h20] = 32'b00000000000000000000000000000000;
assign rom[6'h21] = 32'b00000000000000000000000000000000;
assign rom[6'h22] = 32'b00000000000000000000000000000000;
assign rom[6'h23] = 32'b00000000000000000000000000000000;
assign rom[6'h24] = 32'b00000000000000000000000000000000;
assign rom[6'h25] = 32'b00000000000000000000000000000000;
assign rom[6'h26] = 32'b00000000000000000000000000000000;
assign rom[6'h27] = 32'b00000000000000000000000000000000;
assign rom[6'h28] = 32'b00000000000000000000000000000000;
assign rom[6'h29] = 32'b00000000000000000000000000000000;
assign rom[6'h2a] = 32'b00000000000000000000000000000000;
assign rom[6'h2b] = 32'b00000000000000000000000000000000;
assign rom[6'h2c] = 32'b00000000000000000000000000000000;
assign rom[6'h2d] = 32'b00000000000000000000000000000000;
assign rom[6'h2e] = 32'b00000000000000000000000000000000;
assign rom[6'h2f] = 32'b00000000000000000000000000000000;
assign rom[6'h30] = 32'b00000000000000000000000000000000;
assign rom[6'h31] = 32'b00000000000000000000000000000000;
assign rom[6'h32] = 32'b00000000000000000000000000000000;
assign rom[6'h33] = 32'b00000000000000000000000000000000;
assign rom[6'h34] = 32'b00000000000000000000000000000000;
assign rom[6'h35] = 32'b00000000000000000000000000000000;
assign rom[6'h36] = 32'b00000000000000000000000000000000;
assign rom[6'h37] = 32'b00000000000000000000000000000000;
assign rom[6'h38] = 32'b00000000000000000000000000000000;
assign rom[6'h39] = 32'b00000000000000000000000000000000;
assign rom[6'h3a] = 32'b00000000000000000000000000000000;
assign rom[6'h3b] = 32'b00000000000000000000000000000000;
assign rom[6'h3c] = 32'b00000000000000000000000000000000;
assign rom[6'h3d] = 32'b00000000000000000000000000000000;
assign rom[6'h3e] = 32'b00000000000000000000000000000000;
assign rom[6'h3f] = 32'b00000000000000000000000000000000;
endmodule
