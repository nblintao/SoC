module inst_mem_v (clk,a,inst,ram_a,d_f_ram,wram,d_t_ram,led_num);
    input clk;
    input  [31:0] a;
    output [31:0] inst; 
    input  [31:0] ram_a;
    output [31:0] d_f_ram;
    input         wram;
    input  [31:0] d_t_ram;
    output reg [7:0] led_num;

    initial led_num = 0;

    reg   [31:0] ram [0:63];
    assign inst = ram[a[7:2]];
    assign d_f_ram = ram[ram_a[7:2]];

    always @(posedge clk)begin
        if(wram)begin
            led_num = led_num + 1;
            ram[ram_a[7:2]] <= d_t_ram;
        end
    end

    initial begin
        ram[6'h00] = 32'b00000000000000000000000000000000;
        ram[6'h01] = 32'b00000000000000000000000000000000;
        ram[6'h02] = 32'b00000000000000000000000000000000;
        ram[6'h03] = 32'b00100000000000110000000000000000;
        ram[6'h04] = 32'b00100000000101000000000000111110;
        ram[6'h05] = 32'b10101100011101000000000000000000;
        ram[6'h06] = 32'b00111100000000111100000000000000;
        ram[6'h07] = 32'b00100000000101000000000000000000;
        ram[6'h08] = 32'b10001110100100100000000000000000;
        ram[6'h09] = 32'b00001100000000000000000000001110;
        ram[6'h0a] = 32'b00100010100101000000000000000100;
        ram[6'h0b] = 32'b00101010100101010000000010000000;
        ram[6'h0c] = 32'b00010110101000001111111111111011;
        ram[6'h0d] = 32'b00001000000000000000000000100101;
        ram[6'h0e] = 32'b00000011111000001001100000100000;
        ram[6'h0f] = 32'b00100000000010000000000000100000;
        ram[6'h10] = 32'b00100001000010001111111111111100;
        ram[6'h11] = 32'b00000001000100100010100000000110;
        ram[6'h12] = 32'b00001100000000000000000000011000;
        ram[6'h13] = 32'b00101001000010010000000000000100;
        ram[6'h14] = 32'b00010001001000001111111111111011;
        ram[6'h15] = 32'b00100000000001010000000000100000;
        ram[6'h16] = 32'b00001100000000000000000000100010;
        ram[6'h17] = 32'b00000010011000000000000000001000;
        ram[6'h18] = 32'b00110000101001010000000000001111;
        ram[6'h19] = 32'b00100000101001111111111111110110;
        ram[6'h1a] = 32'b00000000000001110011111111000010;
        ram[6'h1b] = 32'b00010000111000000000000000000010;
        ram[6'h1c] = 32'b00100000101001010000000000110000;
        ram[6'h1d] = 32'b00001000000000000000000000011111;
        ram[6'h1e] = 32'b00100000101001010000000000110111;
        ram[6'h1f] = 32'b10101100011001010000000000000000;
        ram[6'h20] = 32'b00100000011000110000000000000100;
        ram[6'h21] = 32'b00000011111000000000000000001000;
        ram[6'h22] = 32'b10101100011001010000000000000000;
        ram[6'h23] = 32'b00100000011000110000000000000100;
        ram[6'h24] = 32'b00000011111000000000000000001000;
        ram[6'h25] = 32'b00001000000000000000000000100101;
        ram[6'h26] = 32'b00000000000000000000000000000000;
        ram[6'h27] = 32'b00000000000000000000000000000000;
        ram[6'h28] = 32'b00000000000000000000000000000000;
        ram[6'h29] = 32'b00000000000000000000000000000000;
        ram[6'h2a] = 32'b00000000000000000000000000000000;
        ram[6'h2b] = 32'b00000000000000000000000000000000;
        ram[6'h2c] = 32'b00000000000000000000000000000000;
        ram[6'h2d] = 32'b00000000000000000000000000000000;
        ram[6'h2e] = 32'b00000000000000000000000000000000;
        ram[6'h2f] = 32'b00000000000000000000000000000000;
        ram[6'h30] = 32'b00000000000000000000000000000000;
        ram[6'h31] = 32'b00000000000000000000000000000000;
        ram[6'h32] = 32'b00000000000000000000000000000000;
        ram[6'h33] = 32'b00000000000000000000000000000000;
        ram[6'h34] = 32'b00000000000000000000000000000000;
        ram[6'h35] = 32'b00000000000000000000000000000000;
        ram[6'h36] = 32'b00000000000000000000000000000000;
        ram[6'h37] = 32'b00000000000000000000000000000000;
        ram[6'h38] = 32'b00000000000000000000000000000000;
        ram[6'h39] = 32'b00000000000000000000000000000000;
        ram[6'h3a] = 32'b00000000000000000000000000000000;
        ram[6'h3b] = 32'b00000000000000000000000000000000;
        ram[6'h3c] = 32'b00000000000000000000000000000000;
        ram[6'h3d] = 32'b00000000000000000000000000000000;
        ram[6'h3e] = 32'b00000000000000000000000000000000;
        ram[6'h3f] = 32'b00000000000000000000000000000000;
    end
endmodule
