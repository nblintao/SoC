`timescale 1ns / 1ps
// data length is 512
// ram depth is 9
module mio_rom (a, inst, rom_a, d_f_rom);
    input  [31:0] a;
    output [31:0] inst; 
    input  [31:0] rom_a;
    output [31:0] d_f_rom;

    wire   [31:0] rom [0:511];
    assign inst    = rom[a[10:2]];
    assign d_f_rom = rom[rom_a[10:2]];

    assign rom[9'h000] = 32'b00100000000111010001000000000000;
    assign rom[9'h001] = 32'b00100011101111011111111111111000;
    assign rom[9'h002] = 32'b00100000000010000000000000011110;
    assign rom[9'h003] = 32'b10101111101010000000000000000000;
    assign rom[9'h004] = 32'b00100000000010000000000000110001;
    assign rom[9'h005] = 32'b10101111101010000000000000000100;
    assign rom[9'h006] = 32'b00000000000111010010000000100000;
    assign rom[9'h007] = 32'b00001100000000000000000100000110;
    assign rom[9'h008] = 32'b00100011101111011111111111100000;
    assign rom[9'h009] = 32'b10101111101000000000000000000000;
    assign rom[9'h00a] = 32'b10101111101000000000000000000100;
    assign rom[9'h00b] = 32'b00100000000010000000000000000101;
    assign rom[9'h00c] = 32'b10101111101010000000000000001000;
    assign rom[9'h00d] = 32'b10101111101010000000000000001100;
    assign rom[9'h00e] = 32'b10101111101000000000000000010000;
    assign rom[9'h00f] = 32'b00100000000010000000000000000010;
    assign rom[9'h010] = 32'b10101111101010000000000000010100;
    assign rom[9'h011] = 32'b10101111101010000000000000011000;
    assign rom[9'h012] = 32'b10101111101000000000000000011100;
    assign rom[9'h013] = 32'b00100000000010000000000000011111;
    assign rom[9'h014] = 32'b00111100000010011100000000000000;
    assign rom[9'h015] = 32'b00110101001010010000000000000000;
    assign rom[9'h016] = 32'b10101101001010000000000000000000;
    assign rom[9'h017] = 32'b00100011101111011111111111100000;
    assign rom[9'h018] = 32'b00100000000010000000000000001010;
    assign rom[9'h019] = 32'b10101111101010000000000000000000;
    assign rom[9'h01a] = 32'b10101111101000000000000000000100;
    assign rom[9'h01b] = 32'b00100000000010000000000000000111;
    assign rom[9'h01c] = 32'b10101111101010000000000000001000;
    assign rom[9'h01d] = 32'b10101111101010000000000000001100;
    assign rom[9'h01e] = 32'b10101111101000000000000000010000;
    assign rom[9'h01f] = 32'b00100000000010000000000000000011;
    assign rom[9'h020] = 32'b10101111101010000000000000010100;
    assign rom[9'h021] = 32'b10101111101010000000000000011000;
    assign rom[9'h022] = 32'b10101111101000000000000000011100;
    assign rom[9'h023] = 32'b00100000000010000000000000011111;
    assign rom[9'h024] = 32'b00111100000010011100000000000000;
    assign rom[9'h025] = 32'b00110101001010010000000000000000;
    assign rom[9'h026] = 32'b10101101001010000000000000000000;
    assign rom[9'h027] = 32'b00111100000010001010000000000000;
    assign rom[9'h028] = 32'b00110101000010000000000000000000;
    assign rom[9'h029] = 32'b10001101000100000000000000000000;
    assign rom[9'h02a] = 32'b00110010000010000000000100000000;
    assign rom[9'h02b] = 32'b00010001000000000000000000000011;
    assign rom[9'h02c] = 32'b00000000000100000010000000000000;
    assign rom[9'h02d] = 32'b00100011101001010000000001000000;
    assign rom[9'h02e] = 32'b00001100000000000000000010011111;
    assign rom[9'h02f] = 32'b10001100000010000001000000001000;
    assign rom[9'h030] = 32'b00010001000000000000000000001011;
    assign rom[9'h031] = 32'b10101100000000000001000000001000;
    assign rom[9'h032] = 32'b00100011101001010000000000000000;
    assign rom[9'h033] = 32'b00001100000000000000000000111101;
    assign rom[9'h034] = 32'b00100011101001000000000001000000;
    assign rom[9'h035] = 32'b00100011101001010000000000000000;
    assign rom[9'h036] = 32'b00001100000000000000000001100100;
    assign rom[9'h037] = 32'b00100011101001010000000000100000;
    assign rom[9'h038] = 32'b00001100000000000000000000111101;
    assign rom[9'h039] = 32'b00100011101001000000000001000000;
    assign rom[9'h03a] = 32'b00100011101001010000000000100000;
    assign rom[9'h03b] = 32'b00001100000000000000000001100100;
    assign rom[9'h03c] = 32'b00001000000000000000000000100111;
    assign rom[9'h03d] = 32'b10001100101010000000000000001100;
    assign rom[9'h03e] = 32'b00010001000000000000000000000011;
    assign rom[9'h03f] = 32'b00100001000010001111111111111111;
    assign rom[9'h040] = 32'b10101100101010000000000000001100;
    assign rom[9'h041] = 32'b00000011111000000000000000001000;
    assign rom[9'h042] = 32'b10001100101010000000000000001000;
    assign rom[9'h043] = 32'b10101100101010000000000000001100;
    assign rom[9'h044] = 32'b10001100101010100000000000000000;
    assign rom[9'h045] = 32'b10001100101010110000000000000100;
    assign rom[9'h046] = 32'b10001100101011000000000000010000;
    assign rom[9'h047] = 32'b00100000000010010000000001001111;
    assign rom[9'h048] = 32'b00010101001010110000000000000100;
    assign rom[9'h049] = 32'b00010101100000000000000000000011;
    assign rom[9'h04a] = 32'b00100000000011000000000000000001;
    assign rom[9'h04b] = 32'b10101100101011000000000000010000;
    assign rom[9'h04c] = 32'b00001000000000000000000001100011;
    assign rom[9'h04d] = 32'b00100000000010010000000000000000;
    assign rom[9'h04e] = 32'b00010101001010110000000000000100;
    assign rom[9'h04f] = 32'b00010001100000000000000000000011;
    assign rom[9'h050] = 32'b00100000000011000000000000000000;
    assign rom[9'h051] = 32'b10101100101011000000000000010000;
    assign rom[9'h052] = 32'b00001000000000000000000001100011;
    assign rom[9'h053] = 32'b00100011101111011111111111110100;
    assign rom[9'h054] = 32'b10101111101001000000000000000000;
    assign rom[9'h055] = 32'b10101111101001010000000000000100;
    assign rom[9'h056] = 32'b10101111101111110000000000001000;
    assign rom[9'h057] = 32'b00000000000010100010000000000000;
    assign rom[9'h058] = 32'b00000000000010110010100000000000;
    assign rom[9'h059] = 32'b00010101100000000000000000000010;
    assign rom[9'h05a] = 32'b00001100000000000000000011001010;
    assign rom[9'h05b] = 32'b00001000000000000000000001011101;
    assign rom[9'h05c] = 32'b00001100000000000000000011011001;
    assign rom[9'h05d] = 32'b10001111101001000000000000000000;
    assign rom[9'h05e] = 32'b10001111101001010000000000000100;
    assign rom[9'h05f] = 32'b10001111101111110000000000001000;
    assign rom[9'h060] = 32'b00100011101111010000000000001100;
    assign rom[9'h061] = 32'b10101100101000100000000000000000;
    assign rom[9'h062] = 32'b10101100101000110000000000000100;
    assign rom[9'h063] = 32'b00000011111000000000000000001000;
    assign rom[9'h064] = 32'b10001100101010000000000000011000;
    assign rom[9'h065] = 32'b00010001000000000000000000000011;
    assign rom[9'h066] = 32'b00100001000010001111111111111111;
    assign rom[9'h067] = 32'b10101100101010000000000000011000;
    assign rom[9'h068] = 32'b00000011111000000000000000001000;
    assign rom[9'h069] = 32'b10001100101010000000000000010100;
    assign rom[9'h06a] = 32'b10101100101010000000000000011000;
    assign rom[9'h06b] = 32'b10001100101010100000000000000000;
    assign rom[9'h06c] = 32'b10001100101010110000000000000100;
    assign rom[9'h06d] = 32'b10001100101011000000000000011100;
    assign rom[9'h06e] = 32'b00100000000010010000000000111010;
    assign rom[9'h06f] = 32'b00010101001010100000000000011000;
    assign rom[9'h070] = 32'b00010101100000000000000000010111;
    assign rom[9'h071] = 32'b00100000000011000000000000000001;
    assign rom[9'h072] = 32'b10101100101011000000000000011100;
    assign rom[9'h073] = 32'b10001100100011010000000000000000;
    assign rom[9'h074] = 32'b10001100100011100000000000000100;
    assign rom[9'h075] = 32'b00000001011011010111100000101010;
    assign rom[9'h076] = 32'b00010101111000000000000000000111;
    assign rom[9'h077] = 32'b00000001110010110111100000101010;
    assign rom[9'h078] = 32'b00010101111000000000000000000101;
    assign rom[9'h079] = 32'b00100001101011010000000000000001;
    assign rom[9'h07a] = 32'b10101100100011010000000000000000;
    assign rom[9'h07b] = 32'b00100001110011101111111111111111;
    assign rom[9'h07c] = 32'b10101100100011100000000000000100;
    assign rom[9'h07d] = 32'b00001000000000000000000010000010;
    assign rom[9'h07e] = 32'b00100001101011011111111111111111;
    assign rom[9'h07f] = 32'b10101100100011010000000000000000;
    assign rom[9'h080] = 32'b00100001110011100000000000000001;
    assign rom[9'h081] = 32'b10101100100011100000000000000100;
    assign rom[9'h082] = 32'b00100011101111011111111111111100;
    assign rom[9'h083] = 32'b10101111101111110000000000000000;
    assign rom[9'h084] = 32'b00001100000000000000000100000110;
    assign rom[9'h085] = 32'b10001111101111110000000000000000;
    assign rom[9'h086] = 32'b00100011101111010000000000000100;
    assign rom[9'h087] = 32'b00001000000000000000000010011110;
    assign rom[9'h088] = 32'b00100000000010010000000000000000;
    assign rom[9'h089] = 32'b00010101001010100000000000000100;
    assign rom[9'h08a] = 32'b00010001100000000000000000000011;
    assign rom[9'h08b] = 32'b00100000000011000000000000000000;
    assign rom[9'h08c] = 32'b10101100101011000000000000011100;
    assign rom[9'h08d] = 32'b00001000000000000000000010011110;
    assign rom[9'h08e] = 32'b00100011101111011111111111110100;
    assign rom[9'h08f] = 32'b10101111101001000000000000000000;
    assign rom[9'h090] = 32'b10101111101001010000000000000100;
    assign rom[9'h091] = 32'b10101111101111110000000000001000;
    assign rom[9'h092] = 32'b00000000000010100010000000000000;
    assign rom[9'h093] = 32'b00000000000010110010100000000000;
    assign rom[9'h094] = 32'b00010101100000000000000000000010;
    assign rom[9'h095] = 32'b00001100000000000000000011101000;
    assign rom[9'h096] = 32'b00001000000000000000000010011000;
    assign rom[9'h097] = 32'b00001100000000000000000011110111;
    assign rom[9'h098] = 32'b10001111101001000000000000000000;
    assign rom[9'h099] = 32'b10001111101001010000000000000100;
    assign rom[9'h09a] = 32'b10001111101111110000000000001000;
    assign rom[9'h09b] = 32'b00100011101111010000000000001100;
    assign rom[9'h09c] = 32'b10101100101000100000000000000000;
    assign rom[9'h09d] = 32'b10101100101000110000000000000100;
    assign rom[9'h09e] = 32'b00000011111000000000000000001000;
    assign rom[9'h09f] = 32'b00100011101111011111111111111100;
    assign rom[9'h0a0] = 32'b10101111101111110000000000000000;
    assign rom[9'h0a1] = 32'b00110000100001000000000011111111;
    assign rom[9'h0a2] = 32'b00100000000010100000000001110100;
    assign rom[9'h0a3] = 32'b00010001010001000000000000001110;
    assign rom[9'h0a4] = 32'b00100000000010100000000001101011;
    assign rom[9'h0a5] = 32'b00010001010001000000000000010111;
    assign rom[9'h0a6] = 32'b00100000000010100000000001001101;
    assign rom[9'h0a7] = 32'b00010001010001000000000000000001;
    assign rom[9'h0a8] = 32'b00001000000000000000000011000111;
    assign rom[9'h0a9] = 32'b00111100000010001010000000000000;
    assign rom[9'h0aa] = 32'b00110101000010000000000000000000;
    assign rom[9'h0ab] = 32'b10001101000010010000000000000000;
    assign rom[9'h0ac] = 32'b00110001001010000000000100000000;
    assign rom[9'h0ad] = 32'b00010001000000001111111111111011;
    assign rom[9'h0ae] = 32'b00110001001010010000000011111111;
    assign rom[9'h0af] = 32'b00100000000010100000000000101101;
    assign rom[9'h0b0] = 32'b00010101010010011111111111111000;
    assign rom[9'h0b1] = 32'b00001000000000000000000011000111;
    assign rom[9'h0b2] = 32'b10001100101010000000000000000000;
    assign rom[9'h0b3] = 32'b10001100101010010000000000000100;
    assign rom[9'h0b4] = 32'b00101001001010100000000001001111;
    assign rom[9'h0b5] = 32'b00010001010000000000000000010001;
    assign rom[9'h0b6] = 32'b00100001000010000000000000000001;
    assign rom[9'h0b7] = 32'b00100001001010010000000000000001;
    assign rom[9'h0b8] = 32'b10101100101010000000000000000000;
    assign rom[9'h0b9] = 32'b10101100101010010000000000000100;
    assign rom[9'h0ba] = 32'b00000000000001010010000000100000;
    assign rom[9'h0bb] = 32'b00001100000000000000000100000110;
    assign rom[9'h0bc] = 32'b00001000000000000000000011000111;
    assign rom[9'h0bd] = 32'b10001100101010000000000000000000;
    assign rom[9'h0be] = 32'b10001100101010010000000000000100;
    assign rom[9'h0bf] = 32'b00010001000000000000000000000111;
    assign rom[9'h0c0] = 32'b00100001000010001111111111111111;
    assign rom[9'h0c1] = 32'b00100001001010011111111111111111;
    assign rom[9'h0c2] = 32'b10101100101010000000000000000000;
    assign rom[9'h0c3] = 32'b10101100101010010000000000000100;
    assign rom[9'h0c4] = 32'b00000000000001010010000000100000;
    assign rom[9'h0c5] = 32'b00001100000000000000000100000110;
    assign rom[9'h0c6] = 32'b00001000000000000000000011000111;
    assign rom[9'h0c7] = 32'b10001111101111110000000000000000;
    assign rom[9'h0c8] = 32'b00100011101111010000000000000100;
    assign rom[9'h0c9] = 32'b00000011111000000000000000001000;
    assign rom[9'h0ca] = 32'b00000000000001000100000110000000;
    assign rom[9'h0cb] = 32'b00000000000001000100100100000000;
    assign rom[9'h0cc] = 32'b00000001000010010100000000100000;
    assign rom[9'h0cd] = 32'b00000001000001010100000000100000;
    assign rom[9'h0ce] = 32'b00000000000010000100000010000000;
    assign rom[9'h0cf] = 32'b00111100000010011100000000000000;
    assign rom[9'h0d0] = 32'b00110101001010010000000000000000;
    assign rom[9'h0d1] = 32'b00000001001010000100100000100000;
    assign rom[9'h0d2] = 32'b00100000000010100000000000011111;
    assign rom[9'h0d3] = 32'b10101101001000000000000000000000;
    assign rom[9'h0d4] = 32'b00100000100000100000000000000000;
    assign rom[9'h0d5] = 32'b00100000101000110000000000000001;
    assign rom[9'h0d6] = 32'b00100001001010010000000000000100;
    assign rom[9'h0d7] = 32'b10101101001010100000000000000000;
    assign rom[9'h0d8] = 32'b00000011111000000000000000001000;
    assign rom[9'h0d9] = 32'b00000000000001000100000110000000;
    assign rom[9'h0da] = 32'b00000000000001000100100100000000;
    assign rom[9'h0db] = 32'b00000001000010010100000000100000;
    assign rom[9'h0dc] = 32'b00000001000001010100000000100000;
    assign rom[9'h0dd] = 32'b00000000000010000100000010000000;
    assign rom[9'h0de] = 32'b00111100000010011100000000000000;
    assign rom[9'h0df] = 32'b00110101001010010000000000000000;
    assign rom[9'h0e0] = 32'b00000001001010000100100000100000;
    assign rom[9'h0e1] = 32'b00100000000010100000000000011111;
    assign rom[9'h0e2] = 32'b10101101001000000000000000000000;
    assign rom[9'h0e3] = 32'b00100000100000100000000000000000;
    assign rom[9'h0e4] = 32'b00100000101000111111111111111111;
    assign rom[9'h0e5] = 32'b00100001001010011111111111111100;
    assign rom[9'h0e6] = 32'b10101101001010100000000000000000;
    assign rom[9'h0e7] = 32'b00000011111000000000000000001000;
    assign rom[9'h0e8] = 32'b00000000000001000100000110000000;
    assign rom[9'h0e9] = 32'b00000000000001000100100100000000;
    assign rom[9'h0ea] = 32'b00000001000010010100000000100000;
    assign rom[9'h0eb] = 32'b00000001000001010100000000100000;
    assign rom[9'h0ec] = 32'b00000000000010000100000010000000;
    assign rom[9'h0ed] = 32'b00111100000010011100000000000000;
    assign rom[9'h0ee] = 32'b00110101001010010000000000000000;
    assign rom[9'h0ef] = 32'b00000001001010000100100000100000;
    assign rom[9'h0f0] = 32'b00100000000010100000000000011111;
    assign rom[9'h0f1] = 32'b10101101001000000000000000000000;
    assign rom[9'h0f2] = 32'b00100000100000100000000000000001;
    assign rom[9'h0f3] = 32'b00100000101000110000000000000000;
    assign rom[9'h0f4] = 32'b00100001001010010000000101000000;
    assign rom[9'h0f5] = 32'b10101101001010100000000000000000;
    assign rom[9'h0f6] = 32'b00000011111000000000000000001000;
    assign rom[9'h0f7] = 32'b00000000000001000100000110000000;
    assign rom[9'h0f8] = 32'b00000000000001000100100100000000;
    assign rom[9'h0f9] = 32'b00000001000010010100000000100000;
    assign rom[9'h0fa] = 32'b00000001000001010100000000100000;
    assign rom[9'h0fb] = 32'b00000000000010000100000010000000;
    assign rom[9'h0fc] = 32'b00111100000010011100000000000000;
    assign rom[9'h0fd] = 32'b00110101001010010000000000000000;
    assign rom[9'h0fe] = 32'b00000001001010000100100000100000;
    assign rom[9'h0ff] = 32'b00100000000010100000000000011111;
    assign rom[9'h100] = 32'b10101101001000000000000000000000;
    assign rom[9'h101] = 32'b00100000100000101111111111111111;
    assign rom[9'h102] = 32'b00100000101000110000000000000000;
    assign rom[9'h103] = 32'b00100001001010011111111011000000;
    assign rom[9'h104] = 32'b10101101001010100000000000000000;
    assign rom[9'h105] = 32'b00000011111000000000000000001000;
    assign rom[9'h106] = 32'b10001100100010000000000000000000;
    assign rom[9'h107] = 32'b10001100100010010000000000000100;
    assign rom[9'h108] = 32'b00111100000010101100000000000000;
    assign rom[9'h109] = 32'b00110101010010100000000000000000;
    assign rom[9'h10a] = 32'b00100001010010100100100111000000;
    assign rom[9'h10b] = 32'b00100001010010110000000101000000;
    assign rom[9'h10c] = 32'b00000000000010000100000010000000;
    assign rom[9'h10d] = 32'b00000000000010010100100010000000;
    assign rom[9'h10e] = 32'b00000001000010100100000000100000;
    assign rom[9'h10f] = 32'b00000001001010100100100000100000;
    assign rom[9'h110] = 32'b00000001010010000110000000101010;
    assign rom[9'h111] = 32'b00010001100000000000000000000010;
    assign rom[9'h112] = 32'b10101101010000000000000000000000;
    assign rom[9'h113] = 32'b00001000000000000000000100011100;
    assign rom[9'h114] = 32'b00000001001010100110000000101010;
    assign rom[9'h115] = 32'b00010101100000000000000000000011;
    assign rom[9'h116] = 32'b00100000000011000000000001111111;
    assign rom[9'h117] = 32'b10101101010011000000000000000000;
    assign rom[9'h118] = 32'b00001000000000000000000100011100;
    assign rom[9'h119] = 32'b00000001010010110110000000101010;
    assign rom[9'h11a] = 32'b00010001100000000000000000000011;
    assign rom[9'h11b] = 32'b10101101010000000000000000000000;
    assign rom[9'h11c] = 32'b00100001010010100000000000000100;
    assign rom[9'h11d] = 32'b00001000000000000000000100010000;
    assign rom[9'h11e] = 32'b00000011111000000000000000001000;
    assign rom[9'h11f] = 32'b00001000000000000000000100011111;
    assign rom[9'h120] = 32'b00000000000000000000000000000000;
    assign rom[9'h121] = 32'b00000000000000000000000000000000;
    assign rom[9'h122] = 32'b00000000000000000000000000000000;
    assign rom[9'h123] = 32'b00000000000000000000000000000000;
    assign rom[9'h124] = 32'b00000000000000000000000000000000;
    assign rom[9'h125] = 32'b00000000000000000000000000000000;
    assign rom[9'h126] = 32'b00000000000000000000000000000000;
    assign rom[9'h127] = 32'b00000000000000000000000000000000;
    assign rom[9'h128] = 32'b00000000000000000000000000000000;
    assign rom[9'h129] = 32'b00000000000000000000000000000000;
    assign rom[9'h12a] = 32'b00000000000000000000000000000000;
    assign rom[9'h12b] = 32'b00000000000000000000000000000000;
    assign rom[9'h12c] = 32'b00000000000000000000000000000000;
    assign rom[9'h12d] = 32'b00000000000000000000000000000000;
    assign rom[9'h12e] = 32'b00000000000000000000000000000000;
    assign rom[9'h12f] = 32'b00000000000000000000000000000000;
    assign rom[9'h130] = 32'b00000000000000000000000000000000;
    assign rom[9'h131] = 32'b00000000000000000000000000000000;
    assign rom[9'h132] = 32'b00000000000000000000000000000000;
    assign rom[9'h133] = 32'b00000000000000000000000000000000;
    assign rom[9'h134] = 32'b00000000000000000000000000000000;
    assign rom[9'h135] = 32'b00000000000000000000000000000000;
    assign rom[9'h136] = 32'b00000000000000000000000000000000;
    assign rom[9'h137] = 32'b00000000000000000000000000000000;
    assign rom[9'h138] = 32'b00000000000000000000000000000000;
    assign rom[9'h139] = 32'b00000000000000000000000000000000;
    assign rom[9'h13a] = 32'b00000000000000000000000000000000;
    assign rom[9'h13b] = 32'b00000000000000000000000000000000;
    assign rom[9'h13c] = 32'b00000000000000000000000000000000;
    assign rom[9'h13d] = 32'b00000000000000000000000000000000;
    assign rom[9'h13e] = 32'b00000000000000000000000000000000;
    assign rom[9'h13f] = 32'b00000000000000000000000000000000;
    assign rom[9'h140] = 32'b00000000000000000000000000000000;
    assign rom[9'h141] = 32'b00000000000000000000000000000000;
    assign rom[9'h142] = 32'b00000000000000000000000000000000;
    assign rom[9'h143] = 32'b00000000000000000000000000000000;
    assign rom[9'h144] = 32'b00000000000000000000000000000000;
    assign rom[9'h145] = 32'b00000000000000000000000000000000;
    assign rom[9'h146] = 32'b00000000000000000000000000000000;
    assign rom[9'h147] = 32'b00000000000000000000000000000000;
    assign rom[9'h148] = 32'b00000000000000000000000000000000;
    assign rom[9'h149] = 32'b00000000000000000000000000000000;
    assign rom[9'h14a] = 32'b00000000000000000000000000000000;
    assign rom[9'h14b] = 32'b00000000000000000000000000000000;
    assign rom[9'h14c] = 32'b00000000000000000000000000000000;
    assign rom[9'h14d] = 32'b00000000000000000000000000000000;
    assign rom[9'h14e] = 32'b00000000000000000000000000000000;
    assign rom[9'h14f] = 32'b00000000000000000000000000000000;
    assign rom[9'h150] = 32'b00000000000000000000000000000000;
    assign rom[9'h151] = 32'b00000000000000000000000000000000;
    assign rom[9'h152] = 32'b00000000000000000000000000000000;
    assign rom[9'h153] = 32'b00000000000000000000000000000000;
    assign rom[9'h154] = 32'b00000000000000000000000000000000;
    assign rom[9'h155] = 32'b00000000000000000000000000000000;
    assign rom[9'h156] = 32'b00000000000000000000000000000000;
    assign rom[9'h157] = 32'b00000000000000000000000000000000;
    assign rom[9'h158] = 32'b00000000000000000000000000000000;
    assign rom[9'h159] = 32'b00000000000000000000000000000000;
    assign rom[9'h15a] = 32'b00000000000000000000000000000000;
    assign rom[9'h15b] = 32'b00000000000000000000000000000000;
    assign rom[9'h15c] = 32'b00000000000000000000000000000000;
    assign rom[9'h15d] = 32'b00000000000000000000000000000000;
    assign rom[9'h15e] = 32'b00000000000000000000000000000000;
    assign rom[9'h15f] = 32'b00000000000000000000000000000000;
    assign rom[9'h160] = 32'b00000000000000000000000000000000;
    assign rom[9'h161] = 32'b00000000000000000000000000000000;
    assign rom[9'h162] = 32'b00000000000000000000000000000000;
    assign rom[9'h163] = 32'b00000000000000000000000000000000;
    assign rom[9'h164] = 32'b00000000000000000000000000000000;
    assign rom[9'h165] = 32'b00000000000000000000000000000000;
    assign rom[9'h166] = 32'b00000000000000000000000000000000;
    assign rom[9'h167] = 32'b00000000000000000000000000000000;
    assign rom[9'h168] = 32'b00000000000000000000000000000000;
    assign rom[9'h169] = 32'b00000000000000000000000000000000;
    assign rom[9'h16a] = 32'b00000000000000000000000000000000;
    assign rom[9'h16b] = 32'b00000000000000000000000000000000;
    assign rom[9'h16c] = 32'b00000000000000000000000000000000;
    assign rom[9'h16d] = 32'b00000000000000000000000000000000;
    assign rom[9'h16e] = 32'b00000000000000000000000000000000;
    assign rom[9'h16f] = 32'b00000000000000000000000000000000;
    assign rom[9'h170] = 32'b00000000000000000000000000000000;
    assign rom[9'h171] = 32'b00000000000000000000000000000000;
    assign rom[9'h172] = 32'b00000000000000000000000000000000;
    assign rom[9'h173] = 32'b00000000000000000000000000000000;
    assign rom[9'h174] = 32'b00000000000000000000000000000000;
    assign rom[9'h175] = 32'b00000000000000000000000000000000;
    assign rom[9'h176] = 32'b00000000000000000000000000000000;
    assign rom[9'h177] = 32'b00000000000000000000000000000000;
    assign rom[9'h178] = 32'b00000000000000000000000000000000;
    assign rom[9'h179] = 32'b00000000000000000000000000000000;
    assign rom[9'h17a] = 32'b00000000000000000000000000000000;
    assign rom[9'h17b] = 32'b00000000000000000000000000000000;
    assign rom[9'h17c] = 32'b00000000000000000000000000000000;
    assign rom[9'h17d] = 32'b00000000000000000000000000000000;
    assign rom[9'h17e] = 32'b00000000000000000000000000000000;
    assign rom[9'h17f] = 32'b00000000000000000000000000000000;
    assign rom[9'h180] = 32'b00000000000000000000000000000000;
    assign rom[9'h181] = 32'b00000000000000000000000000000000;
    assign rom[9'h182] = 32'b00000000000000000000000000000000;
    assign rom[9'h183] = 32'b00000000000000000000000000000000;
    assign rom[9'h184] = 32'b00000000000000000000000000000000;
    assign rom[9'h185] = 32'b00000000000000000000000000000000;
    assign rom[9'h186] = 32'b00000000000000000000000000000000;
    assign rom[9'h187] = 32'b00000000000000000000000000000000;
    assign rom[9'h188] = 32'b00000000000000000000000000000000;
    assign rom[9'h189] = 32'b00000000000000000000000000000000;
    assign rom[9'h18a] = 32'b00000000000000000000000000000000;
    assign rom[9'h18b] = 32'b00000000000000000000000000000000;
    assign rom[9'h18c] = 32'b00000000000000000000000000000000;
    assign rom[9'h18d] = 32'b00000000000000000000000000000000;
    assign rom[9'h18e] = 32'b00000000000000000000000000000000;
    assign rom[9'h18f] = 32'b00000000000000000000000000000000;
    assign rom[9'h190] = 32'b00000000000000000000000000000000;
    assign rom[9'h191] = 32'b00000000000000000000000000000000;
    assign rom[9'h192] = 32'b00000000000000000000000000000000;
    assign rom[9'h193] = 32'b00000000000000000000000000000000;
    assign rom[9'h194] = 32'b00000000000000000000000000000000;
    assign rom[9'h195] = 32'b00000000000000000000000000000000;
    assign rom[9'h196] = 32'b00000000000000000000000000000000;
    assign rom[9'h197] = 32'b00000000000000000000000000000000;
    assign rom[9'h198] = 32'b00000000000000000000000000000000;
    assign rom[9'h199] = 32'b00000000000000000000000000000000;
    assign rom[9'h19a] = 32'b00000000000000000000000000000000;
    assign rom[9'h19b] = 32'b00000000000000000000000000000000;
    assign rom[9'h19c] = 32'b00000000000000000000000000000000;
    assign rom[9'h19d] = 32'b00000000000000000000000000000000;
    assign rom[9'h19e] = 32'b00000000000000000000000000000000;
    assign rom[9'h19f] = 32'b00000000000000000000000000000000;
    assign rom[9'h1a0] = 32'b00000000000000000000000000000000;
    assign rom[9'h1a1] = 32'b00000000000000000000000000000000;
    assign rom[9'h1a2] = 32'b00000000000000000000000000000000;
    assign rom[9'h1a3] = 32'b00000000000000000000000000000000;
    assign rom[9'h1a4] = 32'b00000000000000000000000000000000;
    assign rom[9'h1a5] = 32'b00000000000000000000000000000000;
    assign rom[9'h1a6] = 32'b00000000000000000000000000000000;
    assign rom[9'h1a7] = 32'b00000000000000000000000000000000;
    assign rom[9'h1a8] = 32'b00000000000000000000000000000000;
    assign rom[9'h1a9] = 32'b00000000000000000000000000000000;
    assign rom[9'h1aa] = 32'b00000000000000000000000000000000;
    assign rom[9'h1ab] = 32'b00000000000000000000000000000000;
    assign rom[9'h1ac] = 32'b00000000000000000000000000000000;
    assign rom[9'h1ad] = 32'b00000000000000000000000000000000;
    assign rom[9'h1ae] = 32'b00000000000000000000000000000000;
    assign rom[9'h1af] = 32'b00000000000000000000000000000000;
    assign rom[9'h1b0] = 32'b00000000000000000000000000000000;
    assign rom[9'h1b1] = 32'b00000000000000000000000000000000;
    assign rom[9'h1b2] = 32'b00000000000000000000000000000000;
    assign rom[9'h1b3] = 32'b00000000000000000000000000000000;
    assign rom[9'h1b4] = 32'b00000000000000000000000000000000;
    assign rom[9'h1b5] = 32'b00000000000000000000000000000000;
    assign rom[9'h1b6] = 32'b00000000000000000000000000000000;
    assign rom[9'h1b7] = 32'b00000000000000000000000000000000;
    assign rom[9'h1b8] = 32'b00000000000000000000000000000000;
    assign rom[9'h1b9] = 32'b00000000000000000000000000000000;
    assign rom[9'h1ba] = 32'b00000000000000000000000000000000;
    assign rom[9'h1bb] = 32'b00000000000000000000000000000000;
    assign rom[9'h1bc] = 32'b00000000000000000000000000000000;
    assign rom[9'h1bd] = 32'b00000000000000000000000000000000;
    assign rom[9'h1be] = 32'b00000000000000000000000000000000;
    assign rom[9'h1bf] = 32'b00000000000000000000000000000000;
    assign rom[9'h1c0] = 32'b00000000000000000000000000000000;
    assign rom[9'h1c1] = 32'b00000000000000000000000000000000;
    assign rom[9'h1c2] = 32'b00000000000000000000000000000000;
    assign rom[9'h1c3] = 32'b00000000000000000000000000000000;
    assign rom[9'h1c4] = 32'b00000000000000000000000000000000;
    assign rom[9'h1c5] = 32'b00000000000000000000000000000000;
    assign rom[9'h1c6] = 32'b00000000000000000000000000000000;
    assign rom[9'h1c7] = 32'b00000000000000000000000000000000;
    assign rom[9'h1c8] = 32'b00000000000000000000000000000000;
    assign rom[9'h1c9] = 32'b00000000000000000000000000000000;
    assign rom[9'h1ca] = 32'b00000000000000000000000000000000;
    assign rom[9'h1cb] = 32'b00000000000000000000000000000000;
    assign rom[9'h1cc] = 32'b00000000000000000000000000000000;
    assign rom[9'h1cd] = 32'b00000000000000000000000000000000;
    assign rom[9'h1ce] = 32'b00000000000000000000000000000000;
    assign rom[9'h1cf] = 32'b00000000000000000000000000000000;
    assign rom[9'h1d0] = 32'b00000000000000000000000000000000;
    assign rom[9'h1d1] = 32'b00000000000000000000000000000000;
    assign rom[9'h1d2] = 32'b00000000000000000000000000000000;
    assign rom[9'h1d3] = 32'b00000000000000000000000000000000;
    assign rom[9'h1d4] = 32'b00000000000000000000000000000000;
    assign rom[9'h1d5] = 32'b00000000000000000000000000000000;
    assign rom[9'h1d6] = 32'b00000000000000000000000000000000;
    assign rom[9'h1d7] = 32'b00000000000000000000000000000000;
    assign rom[9'h1d8] = 32'b00000000000000000000000000000000;
    assign rom[9'h1d9] = 32'b00000000000000000000000000000000;
    assign rom[9'h1da] = 32'b00000000000000000000000000000000;
    assign rom[9'h1db] = 32'b00000000000000000000000000000000;
    assign rom[9'h1dc] = 32'b00000000000000000000000000000000;
    assign rom[9'h1dd] = 32'b00000000000000000000000000000000;
    assign rom[9'h1de] = 32'b00000000000000000000000000000000;
    assign rom[9'h1df] = 32'b00000000000000000000000000000000;
    assign rom[9'h1e0] = 32'b00000000000000000000000000000000;
    assign rom[9'h1e1] = 32'b00000000000000000000000000000000;
    assign rom[9'h1e2] = 32'b00000000000000000000000000000000;
    assign rom[9'h1e3] = 32'b00000000000000000000000000000000;
    assign rom[9'h1e4] = 32'b00000000000000000000000000000000;
    assign rom[9'h1e5] = 32'b00000000000000000000000000000000;
    assign rom[9'h1e6] = 32'b00000000000000000000000000000000;
    assign rom[9'h1e7] = 32'b00000000000000000000000000000000;
    assign rom[9'h1e8] = 32'b00000000000000000000000000000000;
    assign rom[9'h1e9] = 32'b00000000000000000000000000000000;
    assign rom[9'h1ea] = 32'b00000000000000000000000000000000;
    assign rom[9'h1eb] = 32'b00000000000000000000000000000000;
    assign rom[9'h1ec] = 32'b00000000000000000000000000000000;
    assign rom[9'h1ed] = 32'b00000000000000000000000000000000;
    assign rom[9'h1ee] = 32'b00000000000000000000000000000000;
    assign rom[9'h1ef] = 32'b00000000000000000000000000000000;
    assign rom[9'h1f0] = 32'b00000000000000000000000000000000;
    assign rom[9'h1f1] = 32'b00000000000000000000000000000000;
    assign rom[9'h1f2] = 32'b00000000000000000000000000000000;
    assign rom[9'h1f3] = 32'b00000000000000000000000000000000;
    assign rom[9'h1f4] = 32'b00000000000000000000000000000000;
    assign rom[9'h1f5] = 32'b00000000000000000000000000000000;
    assign rom[9'h1f6] = 32'b00000000000000000000000000000000;
    assign rom[9'h1f7] = 32'b00000000000000000000000000000000;
    assign rom[9'h1f8] = 32'b00000000000000000000000000000000;
    assign rom[9'h1f9] = 32'b00000000000000000000000000000000;
    assign rom[9'h1fa] = 32'b00000000000000000000000000000000;
    assign rom[9'h1fb] = 32'b00000000000000000000000000000000;
    assign rom[9'h1fc] = 32'b00000000000000000000000000000000;
    assign rom[9'h1fd] = 32'b00000000000000000000000000000000;
    assign rom[9'h1fe] = 32'b00000000000000000000000000000000;
    assign rom[9'h1ff] = 32'b00000000000000000000000000000000;
endmodule
